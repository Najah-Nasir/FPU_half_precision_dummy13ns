##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Tue May 31 00:36:02 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 1020.280000 BY 1019.660000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.852 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8708 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.193 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 144.448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 771.328 LAYER met3  ;
    ANTENNAGATEAREA 0.852 LAYER met3  ;
    ANTENNAMAXAREACAR 170.052 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 906.867 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.107277 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2.015000 0.000000 2.155000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.131 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 57.8188 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 285.061 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 5.200000 0.490000 5.340000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.875000 0.000000 217.015000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.940000 0.000000 73.080000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.960000 0.000000 219.100000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.790000 0.000000 214.930000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.700000 0.000000 212.840000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.615000 0.000000 210.755000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.530000 0.000000 208.670000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.690000 0.000000 139.830000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.605000 0.000000 137.745000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.520000 0.000000 135.660000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.435000 0.000000 133.575000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.350000 0.000000 131.490000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.260000 0.000000 129.400000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.175000 0.000000 127.315000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.090000 0.000000 125.230000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.005000 0.000000 123.145000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.920000 0.000000 121.060000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.830000 0.000000 118.970000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.745000 0.000000 116.885000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.660000 0.000000 114.800000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.575000 0.000000 112.715000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490000 0.000000 110.630000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.400000 0.000000 108.540000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.315000 0.000000 106.455000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.230000 0.000000 104.370000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.145000 0.000000 102.285000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.060000 0.000000 100.200000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.970000 0.000000 98.110000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.885000 0.000000 96.025000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.800000 0.000000 93.940000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.715000 0.000000 91.855000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.630000 0.000000 89.770000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.540000 0.000000 87.680000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.455000 0.000000 85.595000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.370000 0.000000 83.510000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.285000 0.000000 81.425000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.200000 0.000000 79.340000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.110000 0.000000 77.250000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.025000 0.000000 75.165000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.855000 0.000000 70.995000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.770000 0.000000 68.910000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.680000 0.000000 66.820000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.595000 0.000000 64.735000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510000 0.000000 62.650000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.425000 0.000000 60.565000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.340000 0.000000 58.480000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.250000 0.000000 56.390000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.165000 0.000000 54.305000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.080000 0.000000 52.220000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.995000 0.000000 50.135000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.910000 0.000000 48.050000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.820000 0.000000 45.960000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.735000 0.000000 43.875000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.650000 0.000000 41.790000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.565000 0.000000 39.705000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.480000 0.000000 37.620000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.390000 0.000000 35.530000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.305000 0.000000 33.445000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.220000 0.000000 31.360000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.135000 0.000000 29.275000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.050000 0.000000 27.190000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.960000 0.000000 25.100000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.875000 0.000000 23.015000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790000 0.000000 20.930000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.705000 0.000000 18.845000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.620000 0.000000 16.760000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.530000 0.000000 14.670000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.445000 0.000000 12.585000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.360000 0.000000 10.500000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.275000 0.000000 8.415000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.190000 0.000000 6.330000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 4.100000 0.000000 4.240000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 206.445000 0.000000 206.585000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 204.360000 0.000000 204.500000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 202.270000 0.000000 202.410000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 200.185000 0.000000 200.325000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 198.100000 0.000000 198.240000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 196.015000 0.000000 196.155000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 193.930000 0.000000 194.070000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 191.840000 0.000000 191.980000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 189.755000 0.000000 189.895000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 187.670000 0.000000 187.810000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 185.585000 0.000000 185.725000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 183.500000 0.000000 183.640000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 181.410000 0.000000 181.550000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 179.325000 0.000000 179.465000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 177.240000 0.000000 177.380000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 175.155000 0.000000 175.295000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 173.070000 0.000000 173.210000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 170.980000 0.000000 171.120000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 168.895000 0.000000 169.035000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 166.810000 0.000000 166.950000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 164.725000 0.000000 164.865000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 162.640000 0.000000 162.780000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 160.550000 0.000000 160.690000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 158.465000 0.000000 158.605000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 156.380000 0.000000 156.520000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 154.295000 0.000000 154.435000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 152.210000 0.000000 152.350000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 150.120000 0.000000 150.260000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 148.035000 0.000000 148.175000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 145.950000 0.000000 146.090000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 143.865000 0.000000 144.005000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 141.780000 0.000000 141.920000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.970000 0.000000 486.110000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.880000 0.000000 484.020000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.795000 0.000000 481.935000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.710000 0.000000 479.850000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.625000 0.000000 477.765000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.540000 0.000000 475.680000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.450000 0.000000 473.590000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.365000 0.000000 471.505000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.280000 0.000000 469.420000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.195000 0.000000 467.335000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.110000 0.000000 465.250000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.020000 0.000000 463.160000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.935000 0.000000 461.075000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.850000 0.000000 458.990000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.765000 0.000000 456.905000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.680000 0.000000 454.820000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.590000 0.000000 452.730000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.505000 0.000000 450.645000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.420000 0.000000 448.560000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.335000 0.000000 446.475000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.250000 0.000000 444.390000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.160000 0.000000 442.300000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.075000 0.000000 440.215000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.990000 0.000000 438.130000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.905000 0.000000 436.045000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.820000 0.000000 433.960000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.730000 0.000000 431.870000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.645000 0.000000 429.785000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.560000 0.000000 427.700000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.475000 0.000000 425.615000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.390000 0.000000 423.530000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.300000 0.000000 421.440000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.215000 0.000000 419.355000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.130000 0.000000 417.270000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.045000 0.000000 415.185000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.960000 0.000000 413.100000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870000 0.000000 411.010000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.785000 0.000000 408.925000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.700000 0.000000 406.840000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.615000 0.000000 404.755000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.530000 0.000000 402.670000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.440000 0.000000 400.580000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.355000 0.000000 398.495000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.270000 0.000000 396.410000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.185000 0.000000 394.325000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.100000 0.000000 392.240000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.010000 0.000000 390.150000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.925000 0.000000 388.065000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.840000 0.000000 385.980000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.755000 0.000000 383.895000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.670000 0.000000 381.810000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.580000 0.000000 379.720000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.495000 0.000000 377.635000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.410000 0.000000 375.550000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.325000 0.000000 373.465000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.240000 0.000000 371.380000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.150000 0.000000 369.290000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.065000 0.000000 367.205000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.980000 0.000000 365.120000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.895000 0.000000 363.035000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.810000 0.000000 360.950000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.720000 0.000000 358.860000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.96 LAYER met2  ;
    ANTENNAMAXAREACAR 1.32859 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 4.89331 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0259596 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 356.635000 0.000000 356.775000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.7017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.3475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 206.355 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1103.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 11.475 LAYER met4  ;
    ANTENNAMAXAREACAR 88.4287 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 463.724 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.426567 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 354.550000 0.000000 354.690000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.465000 0.000000 352.605000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.380000 0.000000 350.520000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.290000 0.000000 348.430000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.205000 0.000000 346.345000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.120000 0.000000 344.260000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.035000 0.000000 342.175000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.950000 0.000000 340.090000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.860000 0.000000 338.000000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.775000 0.000000 335.915000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.690000 0.000000 333.830000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.605000 0.000000 331.745000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.520000 0.000000 329.660000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.430000 0.000000 327.570000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.345000 0.000000 325.485000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.260000 0.000000 323.400000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.175000 0.000000 321.315000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.090000 0.000000 319.230000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.000000 0.000000 317.140000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.915000 0.000000 315.055000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.830000 0.000000 312.970000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.745000 0.000000 310.885000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.660000 0.000000 308.800000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.570000 0.000000 306.710000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.485000 0.000000 304.625000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.400000 0.000000 302.540000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.315000 0.000000 300.455000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.230000 0.000000 298.370000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.140000 0.000000 296.280000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.055000 0.000000 294.195000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.970000 0.000000 292.110000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.885000 0.000000 290.025000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.800000 0.000000 287.940000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8944 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.364 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.3303 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.2091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.162222 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 285.710000 0.000000 285.850000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.48343 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.1465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 283.625000 0.000000 283.765000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.709 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.81 LAYER met2  ;
    ANTENNAMAXAREACAR 7.97575 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.246 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 281.540000 0.000000 281.680000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 8.78905 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.1611 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 279.455000 0.000000 279.595000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.11 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2375 LAYER met2  ;
    ANTENNAMAXAREACAR 3.99067 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.2823 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 277.370000 0.000000 277.510000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.343 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 18.4274 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.3903 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 275.280000 0.000000 275.420000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2539 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.7958 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 273.195000 0.000000 273.335000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.974 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8255 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.2896 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 271.110000 0.000000 271.250000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5313 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.8271 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 269.025000 0.000000 269.165000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.917 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.45 LAYER met2  ;
    ANTENNAMAXAREACAR 6.274 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.2275 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.192716 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 266.940000 0.000000 267.080000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.61 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 6.60828 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.1455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 264.850000 0.000000 264.990000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8565 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.21879 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.9707 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 262.765000 0.000000 262.905000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3744 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.548 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 10.5291 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.9291 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 260.680000 0.000000 260.820000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 8.26485 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.4737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 258.595000 0.000000 258.735000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.556 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 9.72889 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.6909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.298586 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 256.510000 0.000000 256.650000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.521 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.41508 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.2391 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 254.420000 0.000000 254.560000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.335000 0.000000 252.475000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.250000 0.000000 250.390000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.165000 0.000000 248.305000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.080000 0.000000 246.220000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.990000 0.000000 244.130000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.905000 0.000000 242.045000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.820000 0.000000 239.960000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.735000 0.000000 237.875000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.650000 0.000000 235.790000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.560000 0.000000 233.700000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.475000 0.000000 231.615000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.390000 0.000000 229.530000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.305000 0.000000 227.445000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.220000 0.000000 225.360000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.84 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.8303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 223.130000 0.000000 223.270000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.045000 0.000000 221.185000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 752.975000 0.000000 753.115000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 750.890000 0.000000 751.030000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 748.805000 0.000000 748.945000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 746.720000 0.000000 746.860000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 744.630000 0.000000 744.770000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 742.545000 0.000000 742.685000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 740.460000 0.000000 740.600000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 738.375000 0.000000 738.515000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 736.290000 0.000000 736.430000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 734.200000 0.000000 734.340000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 732.115000 0.000000 732.255000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 730.030000 0.000000 730.170000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 727.945000 0.000000 728.085000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 725.860000 0.000000 726.000000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 723.770000 0.000000 723.910000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 721.685000 0.000000 721.825000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 719.600000 0.000000 719.740000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 717.515000 0.000000 717.655000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 715.430000 0.000000 715.570000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 713.340000 0.000000 713.480000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 711.255000 0.000000 711.395000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 709.170000 0.000000 709.310000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 707.085000 0.000000 707.225000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 705.000000 0.000000 705.140000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 702.910000 0.000000 703.050000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 700.825000 0.000000 700.965000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 698.740000 0.000000 698.880000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 696.655000 0.000000 696.795000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 694.570000 0.000000 694.710000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 692.480000 0.000000 692.620000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 690.395000 0.000000 690.535000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 688.310000 0.000000 688.450000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 686.225000 0.000000 686.365000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 684.140000 0.000000 684.280000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 682.050000 0.000000 682.190000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 679.965000 0.000000 680.105000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 677.880000 0.000000 678.020000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 675.795000 0.000000 675.935000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 673.710000 0.000000 673.850000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 671.620000 0.000000 671.760000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 669.535000 0.000000 669.675000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 667.450000 0.000000 667.590000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 665.365000 0.000000 665.505000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 663.280000 0.000000 663.420000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 661.190000 0.000000 661.330000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 659.105000 0.000000 659.245000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 657.020000 0.000000 657.160000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 654.935000 0.000000 655.075000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 652.850000 0.000000 652.990000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 650.760000 0.000000 650.900000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 648.675000 0.000000 648.815000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 646.590000 0.000000 646.730000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 644.505000 0.000000 644.645000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 642.420000 0.000000 642.560000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 640.330000 0.000000 640.470000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 638.245000 0.000000 638.385000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 636.160000 0.000000 636.300000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 634.075000 0.000000 634.215000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 631.990000 0.000000 632.130000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 629.900000 0.000000 630.040000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 627.815000 0.000000 627.955000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 625.730000 0.000000 625.870000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 623.645000 0.000000 623.785000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 621.560000 0.000000 621.700000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 619.470000 0.000000 619.610000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 617.385000 0.000000 617.525000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 615.300000 0.000000 615.440000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 613.215000 0.000000 613.355000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 611.130000 0.000000 611.270000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 609.040000 0.000000 609.180000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 606.955000 0.000000 607.095000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 604.870000 0.000000 605.010000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 602.785000 0.000000 602.925000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 600.700000 0.000000 600.840000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 598.610000 0.000000 598.750000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 596.525000 0.000000 596.665000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 594.440000 0.000000 594.580000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 592.355000 0.000000 592.495000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 590.270000 0.000000 590.410000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 588.180000 0.000000 588.320000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.122 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.9788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 459.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 586.095000 0.000000 586.235000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.3575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.8588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 458.384 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 584.010000 0.000000 584.150000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.5888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 456.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 581.925000 0.000000 582.065000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 82.7958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 442.048 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 579.840000 0.000000 579.980000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.8789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.1468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 411.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 577.750000 0.000000 577.890000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.02 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.1598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 422.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 575.665000 0.000000 575.805000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.1175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 76.3428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 407.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 573.580000 0.000000 573.720000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.583 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 419.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 571.495000 0.000000 571.635000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.1835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.2538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 369.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 569.410000 0.000000 569.550000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8783 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 77.5518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 414.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 567.320000 0.000000 567.460000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.249 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 71.4018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 381.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 565.235000 0.000000 565.375000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.0345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 74.2818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 396.64 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 563.150000 0.000000 563.290000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.266 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 72.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 389.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 561.065000 0.000000 561.205000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0637 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.1575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.4738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 365.664 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 558.980000 0.000000 559.120000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.0575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 73.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 391.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 556.890000 0.000000 557.030000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7628 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.653 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 76.0878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 406.272 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 554.805000 0.000000 554.945000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 552.720000 0.000000 552.860000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 550.635000 0.000000 550.775000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 548.550000 0.000000 548.690000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 546.460000 0.000000 546.600000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 544.375000 0.000000 544.515000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 542.290000 0.000000 542.430000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 540.205000 0.000000 540.345000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 538.120000 0.000000 538.260000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 536.030000 0.000000 536.170000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 533.945000 0.000000 534.085000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 531.860000 0.000000 532.000000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 529.775000 0.000000 529.915000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 527.690000 0.000000 527.830000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 525.600000 0.000000 525.740000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 523.515000 0.000000 523.655000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 521.430000 0.000000 521.570000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 519.345000 0.000000 519.485000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 517.260000 0.000000 517.400000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 515.170000 0.000000 515.310000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 513.085000 0.000000 513.225000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 511.000000 0.000000 511.140000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 508.915000 0.000000 509.055000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 506.830000 0.000000 506.970000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 504.740000 0.000000 504.880000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 502.655000 0.000000 502.795000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 500.570000 0.000000 500.710000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 498.485000 0.000000 498.625000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 496.400000 0.000000 496.540000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 494.310000 0.000000 494.450000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.773 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 492.225000 0.000000 492.365000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.822 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 490.140000 0.000000 490.280000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.0607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 321.626 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 488.055000 0.000000 488.195000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.920000 0.000000 1015.060000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.900000 0.000000 1018.040000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.810000 0.000000 1015.950000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.725000 0.000000 1013.865000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.640000 0.000000 1011.780000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.555000 0.000000 1009.695000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.470000 0.000000 1007.610000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.380000 0.000000 1005.520000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.295000 0.000000 1003.435000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.210000 0.000000 1001.350000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.125000 0.000000 999.265000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.040000 0.000000 997.180000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.950000 0.000000 995.090000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.865000 0.000000 993.005000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.780000 0.000000 990.920000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.695000 0.000000 988.835000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.610000 0.000000 986.750000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.520000 0.000000 984.660000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.435000 0.000000 982.575000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350000 0.000000 980.490000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.265000 0.000000 978.405000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.180000 0.000000 976.320000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.090000 0.000000 974.230000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.005000 0.000000 972.145000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.920000 0.000000 970.060000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.835000 0.000000 967.975000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.750000 0.000000 965.890000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.660000 0.000000 963.800000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.575000 0.000000 961.715000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.490000 0.000000 959.630000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.405000 0.000000 957.545000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.320000 0.000000 955.460000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.230000 0.000000 953.370000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.145000 0.000000 951.285000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.060000 0.000000 949.200000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.975000 0.000000 947.115000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.890000 0.000000 945.030000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.800000 0.000000 942.940000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.715000 0.000000 940.855000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.630000 0.000000 938.770000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.545000 0.000000 936.685000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.460000 0.000000 934.600000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370000 0.000000 932.510000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.285000 0.000000 930.425000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.200000 0.000000 928.340000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.115000 0.000000 926.255000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.030000 0.000000 924.170000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.940000 0.000000 922.080000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.855000 0.000000 919.995000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.770000 0.000000 917.910000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.685000 0.000000 915.825000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.600000 0.000000 913.740000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.510000 0.000000 911.650000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.425000 0.000000 909.565000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.340000 0.000000 907.480000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.255000 0.000000 905.395000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.170000 0.000000 903.310000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.080000 0.000000 901.220000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.995000 0.000000 899.135000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.910000 0.000000 897.050000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.825000 0.000000 894.965000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.740000 0.000000 892.880000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.612 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.578 LAYER met2  ;
    ANTENNAMAXAREACAR 3.35589 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.8286 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 890.650000 0.000000 890.790000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 223.069 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 172.376 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 921.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.395 LAYER met3  ;
    ANTENNAMAXAREACAR 29.9588 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.548 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.218932 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 137.531 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 735.84 LAYER met4  ;
    ANTENNAGATEAREA 17.3265 LAYER met4  ;
    ANTENNAMAXAREACAR 50.9045 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 254.911 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.334731 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 888.565000 0.000000 888.705000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.480000 0.000000 886.620000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.395000 0.000000 884.535000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.310000 0.000000 882.450000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.220000 0.000000 880.360000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.135000 0.000000 878.275000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.050000 0.000000 876.190000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.965000 0.000000 874.105000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.880000 0.000000 872.020000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.790000 0.000000 869.930000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.705000 0.000000 867.845000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.620000 0.000000 865.760000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.535000 0.000000 863.675000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.450000 0.000000 861.590000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.360000 0.000000 859.500000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.275000 0.000000 857.415000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.190000 0.000000 855.330000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.588 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.88162 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.1455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 853.105000 0.000000 853.245000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.66343 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.5535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 851.020000 0.000000 851.160000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.13778 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.7414 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 848.930000 0.000000 849.070000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2344 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.0061 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 846.845000 0.000000 846.985000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.427 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.6695 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.6293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 844.760000 0.000000 844.900000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2425 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.94727 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0768 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 842.675000 0.000000 842.815000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.427 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.57465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.4939 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 840.590000 0.000000 840.730000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3705 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.87747 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.0687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 838.500000 0.000000 838.640000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.12606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.3677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 836.415000 0.000000 836.555000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.197 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.67394 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.3333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 834.330000 0.000000 834.470000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.40646 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.0849 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 832.245000 0.000000 832.385000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.00414 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.8545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 830.160000 0.000000 830.300000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.30869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.2808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 828.070000 0.000000 828.210000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.85657 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.2465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 825.985000 0.000000 826.125000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.55253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.6101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 823.900000 0.000000 824.040000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.75646 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.6162 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 821.815000 0.000000 821.955000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.739 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.3 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.5263 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 819.730000 0.000000 819.870000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 3.96222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.8374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 817.640000 0.000000 817.780000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9555 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER met2  ;
    ANTENNAMAXAREACAR 3.48767 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.3524 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0892361 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 815.555000 0.000000 815.695000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.16525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.9889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 813.470000 0.000000 813.610000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.304 LAYER met2  ;
    ANTENNAMAXAREACAR 1.74763 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 6.65148 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.022309 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 811.385000 0.000000 811.525000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 1.91569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.73655 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 809.300000 0.000000 809.440000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.961 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.99051 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.8596 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 807.210000 0.000000 807.350000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.70626 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.8162 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 805.125000 0.000000 805.265000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.76 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.152 LAYER met2  ;
    ANTENNAMAXAREACAR 2.59868 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.1515 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0446181 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 803.040000 0.000000 803.180000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER met2  ;
    ANTENNAMAXAREACAR 3.73715 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.4826 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0892361 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 800.955000 0.000000 801.095000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6778 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.281 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.45717 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.1929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 798.870000 0.000000 799.010000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.861 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.79535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.2616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 796.780000 0.000000 796.920000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.34384 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.7455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 794.695000 0.000000 794.835000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.07253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.3889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 792.610000 0.000000 792.750000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9795 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 6.88485 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.5596 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 790.525000 0.000000 790.665000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.826 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.19414 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.997 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 788.440000 0.000000 788.580000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.350000 0.000000 786.490000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.265000 0.000000 784.405000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.180000 0.000000 782.320000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.095000 0.000000 780.235000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.010000 0.000000 778.150000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.920000 0.000000 776.060000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.835000 0.000000 773.975000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.750000 0.000000 771.890000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.665000 0.000000 769.805000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.580000 0.000000 767.720000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.490000 0.000000 765.630000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.405000 0.000000 763.545000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.320000 0.000000 761.460000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.235000 0.000000 759.375000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.432 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 5.94222 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.8071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 757.150000 0.000000 757.290000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.060000 0.000000 755.200000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 49.590000 0.800000 49.890000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 124.195000 0.800000 124.495000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 198.800000 0.800000 199.100000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 273.410000 0.800000 273.710000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 348.015000 0.800000 348.315000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 422.625000 0.800000 422.925000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 497.230000 0.800000 497.530000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 571.835000 0.800000 572.135000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 646.445000 0.800000 646.745000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 721.050000 0.800000 721.350000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 795.660000 0.800000 795.960000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 870.265000 0.800000 870.565000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 944.870000 0.800000 945.170000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1014.550000 0.800000 1014.850000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.410000 1019.170000 78.550000 1019.660000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.135000 1019.170000 196.275000 1019.660000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.860000 1019.170000 314.000000 1019.660000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.580000 1019.170000 431.720000 1019.660000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.305000 1019.170000 549.445000 1019.660000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.025000 1019.170000 667.165000 1019.660000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.750000 1019.170000 784.890000 1019.660000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.475000 1019.170000 902.615000 1019.660000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.380000 1019.170000 1015.520000 1019.660000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 973.160000 1020.280000 973.460000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 903.635000 1020.280000 903.935000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 834.115000 1020.280000 834.415000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 764.590000 1020.280000 764.890000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 695.070000 1020.280000 695.370000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 625.550000 1020.280000 625.850000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 556.025000 1020.280000 556.325000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 486.505000 1020.280000 486.805000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 416.980000 1020.280000 417.280000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 66.556 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.978 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 347.460000 1020.280000 347.760000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 277.940000 1020.280000 278.240000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 208.415000 1020.280000 208.715000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 138.895000 1020.280000 139.195000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 69.370000 1020.280000 69.670000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 4.390000 1020.280000 4.690000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 24.720000 0.800000 25.020000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 99.325000 0.800000 99.625000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 173.935000 0.800000 174.235000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.79 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 21.9911 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 111.556 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 248.540000 0.800000 248.840000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 323.145000 0.800000 323.445000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 397.755000 0.800000 398.055000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 472.360000 0.800000 472.660000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 546.970000 0.800000 547.270000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 621.575000 0.800000 621.875000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 696.180000 0.800000 696.480000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 770.790000 0.800000 771.090000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 845.395000 0.800000 845.695000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 920.005000 0.800000 920.305000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 994.610000 0.800000 994.910000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 68.1175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 340.309 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.44 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.0998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 39.170000 1019.170000 39.310000 1019.660000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 67.7276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 338.359 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.94 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.4288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 156.895000 1019.170000 157.035000 1019.660000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 162.743 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.7 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 260.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 122.825 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 655.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 274.615000 1019.170000 274.755000 1019.660000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.2469 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 196.074 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.063 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 587.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 392.340000 1019.170000 392.480000 1019.660000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.715 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 176.969 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 944.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 510.065000 1019.170000 510.205000 1019.660000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 79.2426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 395.934 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.622 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.0388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.344 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 627.785000 1019.170000 627.925000 1019.660000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 66.4739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 332.09 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.832 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 196.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.2608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 745.510000 1019.170000 745.650000 1019.660000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.751 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.7838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 249.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 863.230000 1019.170000 863.370000 1019.660000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 70.0264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 349.853 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.35 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.1108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 980.955000 1019.170000 981.095000 1019.660000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 127.869 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 682.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.8318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.24 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 996.330000 1020.280000 996.630000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.2074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.9888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.744 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 926.810000 1020.280000 927.110000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 123.603 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 659.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.7118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 857.290000 1020.280000 857.590000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 127.808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 682.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.5878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.272 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 787.765000 1020.280000 788.065000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5909 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.2348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 718.245000 1020.280000 718.545000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.7934 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.0538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 283.424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 648.720000 1020.280000 649.020000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.4418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.16 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 579.200000 1020.280000 579.500000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 509.680000 1020.280000 509.980000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 440.155000 1020.280000 440.455000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 370.635000 1020.280000 370.935000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 301.110000 1020.280000 301.410000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 231.590000 1020.280000 231.890000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 162.070000 1020.280000 162.370000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 92.545000 1020.280000 92.845000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 23.025000 1020.280000 23.325000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.5 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 4.680000 0.000000 4.980000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 74.455000 0.800000 74.755000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.065000 0.800000 149.365000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 223.670000 0.800000 223.970000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 298.280000 0.800000 298.580000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 372.885000 0.800000 373.185000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 447.490000 0.800000 447.790000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 522.100000 0.800000 522.400000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 596.705000 0.800000 597.005000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 671.315000 0.800000 671.615000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 745.920000 0.800000 746.220000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 820.525000 0.800000 820.825000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 895.135000 0.800000 895.435000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 969.740000 0.800000 970.040000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 5.220000 1019.170000 5.360000 1019.660000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 117.655000 1019.170000 117.795000 1019.660000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 235.375000 1019.170000 235.515000 1019.660000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 353.100000 1019.170000 353.240000 1019.660000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.19 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 470.820000 1019.170000 470.960000 1019.660000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 588.545000 1019.170000 588.685000 1019.660000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 706.270000 1019.170000 706.410000 1019.660000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 823.990000 1019.170000 824.130000 1019.660000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.829 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 442.659 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2388.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 941.715000 1019.170000 941.855000 1019.660000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 1013.940000 1020.280000 1014.240000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 949.985000 1020.280000 950.285000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 880.460000 1020.280000 880.760000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 810.940000 1020.280000 811.240000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 741.420000 1020.280000 741.720000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 671.895000 1020.280000 672.195000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 602.375000 1020.280000 602.675000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 532.850000 1020.280000 533.150000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 463.330000 1020.280000 463.630000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 168.9 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 902.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 12.852 LAYER met3  ;
    ANTENNAMAXAREACAR 35.5508 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 177.659 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.368923 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.7008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.464 LAYER met4  ;
    ANTENNAGATEAREA 15.8715 LAYER met4  ;
    ANTENNAMAXAREACAR 38.1782 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 191.738 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 393.810000 1020.280000 394.110000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 324.285000 1020.280000 324.585000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 254.765000 1020.280000 255.065000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 185.240000 1020.280000 185.540000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 115.720000 1020.280000 116.020000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1019.480000 46.200000 1020.280000 46.500000 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.250000 0.800000 20.550000 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2387.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 0.730000 0.800000 1.030000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 442.419 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2386.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 2.63273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 17.8424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 9.880000 0.800000 10.180000 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1016.220000 1.930000 1018.220000 1016.880000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.060000 1.930000 4.060000 1016.880000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 954.385000 559.895000 956.125000 954.675000 ;
      LAYER met4 ;
        RECT 479.065000 559.895000 480.805000 954.675000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1012.220000 5.930000 1014.220000 1012.880000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.060000 5.930000 8.060000 1012.880000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 482.465000 563.295000 484.205000 951.275000 ;
      LAYER met4 ;
        RECT 950.985000 563.295000 952.725000 951.275000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 1020.280000 1019.660000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 1020.280000 1019.660000 ;
    LAYER met2 ;
      RECT 1015.660000 1019.030000 1020.280000 1019.660000 ;
      RECT 981.235000 1019.030000 1015.240000 1019.660000 ;
      RECT 941.995000 1019.030000 980.815000 1019.660000 ;
      RECT 902.755000 1019.030000 941.575000 1019.660000 ;
      RECT 863.510000 1019.030000 902.335000 1019.660000 ;
      RECT 824.270000 1019.030000 863.090000 1019.660000 ;
      RECT 785.030000 1019.030000 823.850000 1019.660000 ;
      RECT 745.790000 1019.030000 784.610000 1019.660000 ;
      RECT 706.550000 1019.030000 745.370000 1019.660000 ;
      RECT 667.305000 1019.030000 706.130000 1019.660000 ;
      RECT 628.065000 1019.030000 666.885000 1019.660000 ;
      RECT 588.825000 1019.030000 627.645000 1019.660000 ;
      RECT 549.585000 1019.030000 588.405000 1019.660000 ;
      RECT 510.345000 1019.030000 549.165000 1019.660000 ;
      RECT 471.100000 1019.030000 509.925000 1019.660000 ;
      RECT 431.860000 1019.030000 470.680000 1019.660000 ;
      RECT 392.620000 1019.030000 431.440000 1019.660000 ;
      RECT 353.380000 1019.030000 392.200000 1019.660000 ;
      RECT 314.140000 1019.030000 352.960000 1019.660000 ;
      RECT 274.895000 1019.030000 313.720000 1019.660000 ;
      RECT 235.655000 1019.030000 274.475000 1019.660000 ;
      RECT 196.415000 1019.030000 235.235000 1019.660000 ;
      RECT 157.175000 1019.030000 195.995000 1019.660000 ;
      RECT 117.935000 1019.030000 156.755000 1019.660000 ;
      RECT 78.690000 1019.030000 117.515000 1019.660000 ;
      RECT 39.450000 1019.030000 78.270000 1019.660000 ;
      RECT 5.500000 1019.030000 39.030000 1019.660000 ;
      RECT 0.000000 1019.030000 5.080000 1019.660000 ;
      RECT 0.000000 5.480000 1020.280000 1019.030000 ;
      RECT 0.630000 5.060000 1020.280000 5.480000 ;
      RECT 0.000000 0.630000 1020.280000 5.060000 ;
      RECT 1018.180000 0.000000 1020.280000 0.630000 ;
      RECT 1016.090000 0.000000 1017.760000 0.630000 ;
      RECT 1015.200000 0.000000 1015.670000 0.630000 ;
      RECT 1014.005000 0.000000 1014.780000 0.630000 ;
      RECT 1011.920000 0.000000 1013.585000 0.630000 ;
      RECT 1009.835000 0.000000 1011.500000 0.630000 ;
      RECT 1007.750000 0.000000 1009.415000 0.630000 ;
      RECT 1005.660000 0.000000 1007.330000 0.630000 ;
      RECT 1003.575000 0.000000 1005.240000 0.630000 ;
      RECT 1001.490000 0.000000 1003.155000 0.630000 ;
      RECT 999.405000 0.000000 1001.070000 0.630000 ;
      RECT 997.320000 0.000000 998.985000 0.630000 ;
      RECT 995.230000 0.000000 996.900000 0.630000 ;
      RECT 993.145000 0.000000 994.810000 0.630000 ;
      RECT 991.060000 0.000000 992.725000 0.630000 ;
      RECT 988.975000 0.000000 990.640000 0.630000 ;
      RECT 986.890000 0.000000 988.555000 0.630000 ;
      RECT 984.800000 0.000000 986.470000 0.630000 ;
      RECT 982.715000 0.000000 984.380000 0.630000 ;
      RECT 980.630000 0.000000 982.295000 0.630000 ;
      RECT 978.545000 0.000000 980.210000 0.630000 ;
      RECT 976.460000 0.000000 978.125000 0.630000 ;
      RECT 974.370000 0.000000 976.040000 0.630000 ;
      RECT 972.285000 0.000000 973.950000 0.630000 ;
      RECT 970.200000 0.000000 971.865000 0.630000 ;
      RECT 968.115000 0.000000 969.780000 0.630000 ;
      RECT 966.030000 0.000000 967.695000 0.630000 ;
      RECT 963.940000 0.000000 965.610000 0.630000 ;
      RECT 961.855000 0.000000 963.520000 0.630000 ;
      RECT 959.770000 0.000000 961.435000 0.630000 ;
      RECT 957.685000 0.000000 959.350000 0.630000 ;
      RECT 955.600000 0.000000 957.265000 0.630000 ;
      RECT 953.510000 0.000000 955.180000 0.630000 ;
      RECT 951.425000 0.000000 953.090000 0.630000 ;
      RECT 949.340000 0.000000 951.005000 0.630000 ;
      RECT 947.255000 0.000000 948.920000 0.630000 ;
      RECT 945.170000 0.000000 946.835000 0.630000 ;
      RECT 943.080000 0.000000 944.750000 0.630000 ;
      RECT 940.995000 0.000000 942.660000 0.630000 ;
      RECT 938.910000 0.000000 940.575000 0.630000 ;
      RECT 936.825000 0.000000 938.490000 0.630000 ;
      RECT 934.740000 0.000000 936.405000 0.630000 ;
      RECT 932.650000 0.000000 934.320000 0.630000 ;
      RECT 930.565000 0.000000 932.230000 0.630000 ;
      RECT 928.480000 0.000000 930.145000 0.630000 ;
      RECT 926.395000 0.000000 928.060000 0.630000 ;
      RECT 924.310000 0.000000 925.975000 0.630000 ;
      RECT 922.220000 0.000000 923.890000 0.630000 ;
      RECT 920.135000 0.000000 921.800000 0.630000 ;
      RECT 918.050000 0.000000 919.715000 0.630000 ;
      RECT 915.965000 0.000000 917.630000 0.630000 ;
      RECT 913.880000 0.000000 915.545000 0.630000 ;
      RECT 911.790000 0.000000 913.460000 0.630000 ;
      RECT 909.705000 0.000000 911.370000 0.630000 ;
      RECT 907.620000 0.000000 909.285000 0.630000 ;
      RECT 905.535000 0.000000 907.200000 0.630000 ;
      RECT 903.450000 0.000000 905.115000 0.630000 ;
      RECT 901.360000 0.000000 903.030000 0.630000 ;
      RECT 899.275000 0.000000 900.940000 0.630000 ;
      RECT 897.190000 0.000000 898.855000 0.630000 ;
      RECT 895.105000 0.000000 896.770000 0.630000 ;
      RECT 893.020000 0.000000 894.685000 0.630000 ;
      RECT 890.930000 0.000000 892.600000 0.630000 ;
      RECT 888.845000 0.000000 890.510000 0.630000 ;
      RECT 886.760000 0.000000 888.425000 0.630000 ;
      RECT 884.675000 0.000000 886.340000 0.630000 ;
      RECT 882.590000 0.000000 884.255000 0.630000 ;
      RECT 880.500000 0.000000 882.170000 0.630000 ;
      RECT 878.415000 0.000000 880.080000 0.630000 ;
      RECT 876.330000 0.000000 877.995000 0.630000 ;
      RECT 874.245000 0.000000 875.910000 0.630000 ;
      RECT 872.160000 0.000000 873.825000 0.630000 ;
      RECT 870.070000 0.000000 871.740000 0.630000 ;
      RECT 867.985000 0.000000 869.650000 0.630000 ;
      RECT 865.900000 0.000000 867.565000 0.630000 ;
      RECT 863.815000 0.000000 865.480000 0.630000 ;
      RECT 861.730000 0.000000 863.395000 0.630000 ;
      RECT 859.640000 0.000000 861.310000 0.630000 ;
      RECT 857.555000 0.000000 859.220000 0.630000 ;
      RECT 855.470000 0.000000 857.135000 0.630000 ;
      RECT 853.385000 0.000000 855.050000 0.630000 ;
      RECT 851.300000 0.000000 852.965000 0.630000 ;
      RECT 849.210000 0.000000 850.880000 0.630000 ;
      RECT 847.125000 0.000000 848.790000 0.630000 ;
      RECT 845.040000 0.000000 846.705000 0.630000 ;
      RECT 842.955000 0.000000 844.620000 0.630000 ;
      RECT 840.870000 0.000000 842.535000 0.630000 ;
      RECT 838.780000 0.000000 840.450000 0.630000 ;
      RECT 836.695000 0.000000 838.360000 0.630000 ;
      RECT 834.610000 0.000000 836.275000 0.630000 ;
      RECT 832.525000 0.000000 834.190000 0.630000 ;
      RECT 830.440000 0.000000 832.105000 0.630000 ;
      RECT 828.350000 0.000000 830.020000 0.630000 ;
      RECT 826.265000 0.000000 827.930000 0.630000 ;
      RECT 824.180000 0.000000 825.845000 0.630000 ;
      RECT 822.095000 0.000000 823.760000 0.630000 ;
      RECT 820.010000 0.000000 821.675000 0.630000 ;
      RECT 817.920000 0.000000 819.590000 0.630000 ;
      RECT 815.835000 0.000000 817.500000 0.630000 ;
      RECT 813.750000 0.000000 815.415000 0.630000 ;
      RECT 811.665000 0.000000 813.330000 0.630000 ;
      RECT 809.580000 0.000000 811.245000 0.630000 ;
      RECT 807.490000 0.000000 809.160000 0.630000 ;
      RECT 805.405000 0.000000 807.070000 0.630000 ;
      RECT 803.320000 0.000000 804.985000 0.630000 ;
      RECT 801.235000 0.000000 802.900000 0.630000 ;
      RECT 799.150000 0.000000 800.815000 0.630000 ;
      RECT 797.060000 0.000000 798.730000 0.630000 ;
      RECT 794.975000 0.000000 796.640000 0.630000 ;
      RECT 792.890000 0.000000 794.555000 0.630000 ;
      RECT 790.805000 0.000000 792.470000 0.630000 ;
      RECT 788.720000 0.000000 790.385000 0.630000 ;
      RECT 786.630000 0.000000 788.300000 0.630000 ;
      RECT 784.545000 0.000000 786.210000 0.630000 ;
      RECT 782.460000 0.000000 784.125000 0.630000 ;
      RECT 780.375000 0.000000 782.040000 0.630000 ;
      RECT 778.290000 0.000000 779.955000 0.630000 ;
      RECT 776.200000 0.000000 777.870000 0.630000 ;
      RECT 774.115000 0.000000 775.780000 0.630000 ;
      RECT 772.030000 0.000000 773.695000 0.630000 ;
      RECT 769.945000 0.000000 771.610000 0.630000 ;
      RECT 767.860000 0.000000 769.525000 0.630000 ;
      RECT 765.770000 0.000000 767.440000 0.630000 ;
      RECT 763.685000 0.000000 765.350000 0.630000 ;
      RECT 761.600000 0.000000 763.265000 0.630000 ;
      RECT 759.515000 0.000000 761.180000 0.630000 ;
      RECT 757.430000 0.000000 759.095000 0.630000 ;
      RECT 755.340000 0.000000 757.010000 0.630000 ;
      RECT 753.255000 0.000000 754.920000 0.630000 ;
      RECT 751.170000 0.000000 752.835000 0.630000 ;
      RECT 749.085000 0.000000 750.750000 0.630000 ;
      RECT 747.000000 0.000000 748.665000 0.630000 ;
      RECT 744.910000 0.000000 746.580000 0.630000 ;
      RECT 742.825000 0.000000 744.490000 0.630000 ;
      RECT 740.740000 0.000000 742.405000 0.630000 ;
      RECT 738.655000 0.000000 740.320000 0.630000 ;
      RECT 736.570000 0.000000 738.235000 0.630000 ;
      RECT 734.480000 0.000000 736.150000 0.630000 ;
      RECT 732.395000 0.000000 734.060000 0.630000 ;
      RECT 730.310000 0.000000 731.975000 0.630000 ;
      RECT 728.225000 0.000000 729.890000 0.630000 ;
      RECT 726.140000 0.000000 727.805000 0.630000 ;
      RECT 724.050000 0.000000 725.720000 0.630000 ;
      RECT 721.965000 0.000000 723.630000 0.630000 ;
      RECT 719.880000 0.000000 721.545000 0.630000 ;
      RECT 717.795000 0.000000 719.460000 0.630000 ;
      RECT 715.710000 0.000000 717.375000 0.630000 ;
      RECT 713.620000 0.000000 715.290000 0.630000 ;
      RECT 711.535000 0.000000 713.200000 0.630000 ;
      RECT 709.450000 0.000000 711.115000 0.630000 ;
      RECT 707.365000 0.000000 709.030000 0.630000 ;
      RECT 705.280000 0.000000 706.945000 0.630000 ;
      RECT 703.190000 0.000000 704.860000 0.630000 ;
      RECT 701.105000 0.000000 702.770000 0.630000 ;
      RECT 699.020000 0.000000 700.685000 0.630000 ;
      RECT 696.935000 0.000000 698.600000 0.630000 ;
      RECT 694.850000 0.000000 696.515000 0.630000 ;
      RECT 692.760000 0.000000 694.430000 0.630000 ;
      RECT 690.675000 0.000000 692.340000 0.630000 ;
      RECT 688.590000 0.000000 690.255000 0.630000 ;
      RECT 686.505000 0.000000 688.170000 0.630000 ;
      RECT 684.420000 0.000000 686.085000 0.630000 ;
      RECT 682.330000 0.000000 684.000000 0.630000 ;
      RECT 680.245000 0.000000 681.910000 0.630000 ;
      RECT 678.160000 0.000000 679.825000 0.630000 ;
      RECT 676.075000 0.000000 677.740000 0.630000 ;
      RECT 673.990000 0.000000 675.655000 0.630000 ;
      RECT 671.900000 0.000000 673.570000 0.630000 ;
      RECT 669.815000 0.000000 671.480000 0.630000 ;
      RECT 667.730000 0.000000 669.395000 0.630000 ;
      RECT 665.645000 0.000000 667.310000 0.630000 ;
      RECT 663.560000 0.000000 665.225000 0.630000 ;
      RECT 661.470000 0.000000 663.140000 0.630000 ;
      RECT 659.385000 0.000000 661.050000 0.630000 ;
      RECT 657.300000 0.000000 658.965000 0.630000 ;
      RECT 655.215000 0.000000 656.880000 0.630000 ;
      RECT 653.130000 0.000000 654.795000 0.630000 ;
      RECT 651.040000 0.000000 652.710000 0.630000 ;
      RECT 648.955000 0.000000 650.620000 0.630000 ;
      RECT 646.870000 0.000000 648.535000 0.630000 ;
      RECT 644.785000 0.000000 646.450000 0.630000 ;
      RECT 642.700000 0.000000 644.365000 0.630000 ;
      RECT 640.610000 0.000000 642.280000 0.630000 ;
      RECT 638.525000 0.000000 640.190000 0.630000 ;
      RECT 636.440000 0.000000 638.105000 0.630000 ;
      RECT 634.355000 0.000000 636.020000 0.630000 ;
      RECT 632.270000 0.000000 633.935000 0.630000 ;
      RECT 630.180000 0.000000 631.850000 0.630000 ;
      RECT 628.095000 0.000000 629.760000 0.630000 ;
      RECT 626.010000 0.000000 627.675000 0.630000 ;
      RECT 623.925000 0.000000 625.590000 0.630000 ;
      RECT 621.840000 0.000000 623.505000 0.630000 ;
      RECT 619.750000 0.000000 621.420000 0.630000 ;
      RECT 617.665000 0.000000 619.330000 0.630000 ;
      RECT 615.580000 0.000000 617.245000 0.630000 ;
      RECT 613.495000 0.000000 615.160000 0.630000 ;
      RECT 611.410000 0.000000 613.075000 0.630000 ;
      RECT 609.320000 0.000000 610.990000 0.630000 ;
      RECT 607.235000 0.000000 608.900000 0.630000 ;
      RECT 605.150000 0.000000 606.815000 0.630000 ;
      RECT 603.065000 0.000000 604.730000 0.630000 ;
      RECT 600.980000 0.000000 602.645000 0.630000 ;
      RECT 598.890000 0.000000 600.560000 0.630000 ;
      RECT 596.805000 0.000000 598.470000 0.630000 ;
      RECT 594.720000 0.000000 596.385000 0.630000 ;
      RECT 592.635000 0.000000 594.300000 0.630000 ;
      RECT 590.550000 0.000000 592.215000 0.630000 ;
      RECT 588.460000 0.000000 590.130000 0.630000 ;
      RECT 586.375000 0.000000 588.040000 0.630000 ;
      RECT 584.290000 0.000000 585.955000 0.630000 ;
      RECT 582.205000 0.000000 583.870000 0.630000 ;
      RECT 580.120000 0.000000 581.785000 0.630000 ;
      RECT 578.030000 0.000000 579.700000 0.630000 ;
      RECT 575.945000 0.000000 577.610000 0.630000 ;
      RECT 573.860000 0.000000 575.525000 0.630000 ;
      RECT 571.775000 0.000000 573.440000 0.630000 ;
      RECT 569.690000 0.000000 571.355000 0.630000 ;
      RECT 567.600000 0.000000 569.270000 0.630000 ;
      RECT 565.515000 0.000000 567.180000 0.630000 ;
      RECT 563.430000 0.000000 565.095000 0.630000 ;
      RECT 561.345000 0.000000 563.010000 0.630000 ;
      RECT 559.260000 0.000000 560.925000 0.630000 ;
      RECT 557.170000 0.000000 558.840000 0.630000 ;
      RECT 555.085000 0.000000 556.750000 0.630000 ;
      RECT 553.000000 0.000000 554.665000 0.630000 ;
      RECT 550.915000 0.000000 552.580000 0.630000 ;
      RECT 548.830000 0.000000 550.495000 0.630000 ;
      RECT 546.740000 0.000000 548.410000 0.630000 ;
      RECT 544.655000 0.000000 546.320000 0.630000 ;
      RECT 542.570000 0.000000 544.235000 0.630000 ;
      RECT 540.485000 0.000000 542.150000 0.630000 ;
      RECT 538.400000 0.000000 540.065000 0.630000 ;
      RECT 536.310000 0.000000 537.980000 0.630000 ;
      RECT 534.225000 0.000000 535.890000 0.630000 ;
      RECT 532.140000 0.000000 533.805000 0.630000 ;
      RECT 530.055000 0.000000 531.720000 0.630000 ;
      RECT 527.970000 0.000000 529.635000 0.630000 ;
      RECT 525.880000 0.000000 527.550000 0.630000 ;
      RECT 523.795000 0.000000 525.460000 0.630000 ;
      RECT 521.710000 0.000000 523.375000 0.630000 ;
      RECT 519.625000 0.000000 521.290000 0.630000 ;
      RECT 517.540000 0.000000 519.205000 0.630000 ;
      RECT 515.450000 0.000000 517.120000 0.630000 ;
      RECT 513.365000 0.000000 515.030000 0.630000 ;
      RECT 511.280000 0.000000 512.945000 0.630000 ;
      RECT 509.195000 0.000000 510.860000 0.630000 ;
      RECT 507.110000 0.000000 508.775000 0.630000 ;
      RECT 505.020000 0.000000 506.690000 0.630000 ;
      RECT 502.935000 0.000000 504.600000 0.630000 ;
      RECT 500.850000 0.000000 502.515000 0.630000 ;
      RECT 498.765000 0.000000 500.430000 0.630000 ;
      RECT 496.680000 0.000000 498.345000 0.630000 ;
      RECT 494.590000 0.000000 496.260000 0.630000 ;
      RECT 492.505000 0.000000 494.170000 0.630000 ;
      RECT 490.420000 0.000000 492.085000 0.630000 ;
      RECT 488.335000 0.000000 490.000000 0.630000 ;
      RECT 486.250000 0.000000 487.915000 0.630000 ;
      RECT 484.160000 0.000000 485.830000 0.630000 ;
      RECT 482.075000 0.000000 483.740000 0.630000 ;
      RECT 479.990000 0.000000 481.655000 0.630000 ;
      RECT 477.905000 0.000000 479.570000 0.630000 ;
      RECT 475.820000 0.000000 477.485000 0.630000 ;
      RECT 473.730000 0.000000 475.400000 0.630000 ;
      RECT 471.645000 0.000000 473.310000 0.630000 ;
      RECT 469.560000 0.000000 471.225000 0.630000 ;
      RECT 467.475000 0.000000 469.140000 0.630000 ;
      RECT 465.390000 0.000000 467.055000 0.630000 ;
      RECT 463.300000 0.000000 464.970000 0.630000 ;
      RECT 461.215000 0.000000 462.880000 0.630000 ;
      RECT 459.130000 0.000000 460.795000 0.630000 ;
      RECT 457.045000 0.000000 458.710000 0.630000 ;
      RECT 454.960000 0.000000 456.625000 0.630000 ;
      RECT 452.870000 0.000000 454.540000 0.630000 ;
      RECT 450.785000 0.000000 452.450000 0.630000 ;
      RECT 448.700000 0.000000 450.365000 0.630000 ;
      RECT 446.615000 0.000000 448.280000 0.630000 ;
      RECT 444.530000 0.000000 446.195000 0.630000 ;
      RECT 442.440000 0.000000 444.110000 0.630000 ;
      RECT 440.355000 0.000000 442.020000 0.630000 ;
      RECT 438.270000 0.000000 439.935000 0.630000 ;
      RECT 436.185000 0.000000 437.850000 0.630000 ;
      RECT 434.100000 0.000000 435.765000 0.630000 ;
      RECT 432.010000 0.000000 433.680000 0.630000 ;
      RECT 429.925000 0.000000 431.590000 0.630000 ;
      RECT 427.840000 0.000000 429.505000 0.630000 ;
      RECT 425.755000 0.000000 427.420000 0.630000 ;
      RECT 423.670000 0.000000 425.335000 0.630000 ;
      RECT 421.580000 0.000000 423.250000 0.630000 ;
      RECT 419.495000 0.000000 421.160000 0.630000 ;
      RECT 417.410000 0.000000 419.075000 0.630000 ;
      RECT 415.325000 0.000000 416.990000 0.630000 ;
      RECT 413.240000 0.000000 414.905000 0.630000 ;
      RECT 411.150000 0.000000 412.820000 0.630000 ;
      RECT 409.065000 0.000000 410.730000 0.630000 ;
      RECT 406.980000 0.000000 408.645000 0.630000 ;
      RECT 404.895000 0.000000 406.560000 0.630000 ;
      RECT 402.810000 0.000000 404.475000 0.630000 ;
      RECT 400.720000 0.000000 402.390000 0.630000 ;
      RECT 398.635000 0.000000 400.300000 0.630000 ;
      RECT 396.550000 0.000000 398.215000 0.630000 ;
      RECT 394.465000 0.000000 396.130000 0.630000 ;
      RECT 392.380000 0.000000 394.045000 0.630000 ;
      RECT 390.290000 0.000000 391.960000 0.630000 ;
      RECT 388.205000 0.000000 389.870000 0.630000 ;
      RECT 386.120000 0.000000 387.785000 0.630000 ;
      RECT 384.035000 0.000000 385.700000 0.630000 ;
      RECT 381.950000 0.000000 383.615000 0.630000 ;
      RECT 379.860000 0.000000 381.530000 0.630000 ;
      RECT 377.775000 0.000000 379.440000 0.630000 ;
      RECT 375.690000 0.000000 377.355000 0.630000 ;
      RECT 373.605000 0.000000 375.270000 0.630000 ;
      RECT 371.520000 0.000000 373.185000 0.630000 ;
      RECT 369.430000 0.000000 371.100000 0.630000 ;
      RECT 367.345000 0.000000 369.010000 0.630000 ;
      RECT 365.260000 0.000000 366.925000 0.630000 ;
      RECT 363.175000 0.000000 364.840000 0.630000 ;
      RECT 361.090000 0.000000 362.755000 0.630000 ;
      RECT 359.000000 0.000000 360.670000 0.630000 ;
      RECT 356.915000 0.000000 358.580000 0.630000 ;
      RECT 354.830000 0.000000 356.495000 0.630000 ;
      RECT 352.745000 0.000000 354.410000 0.630000 ;
      RECT 350.660000 0.000000 352.325000 0.630000 ;
      RECT 348.570000 0.000000 350.240000 0.630000 ;
      RECT 346.485000 0.000000 348.150000 0.630000 ;
      RECT 344.400000 0.000000 346.065000 0.630000 ;
      RECT 342.315000 0.000000 343.980000 0.630000 ;
      RECT 340.230000 0.000000 341.895000 0.630000 ;
      RECT 338.140000 0.000000 339.810000 0.630000 ;
      RECT 336.055000 0.000000 337.720000 0.630000 ;
      RECT 333.970000 0.000000 335.635000 0.630000 ;
      RECT 331.885000 0.000000 333.550000 0.630000 ;
      RECT 329.800000 0.000000 331.465000 0.630000 ;
      RECT 327.710000 0.000000 329.380000 0.630000 ;
      RECT 325.625000 0.000000 327.290000 0.630000 ;
      RECT 323.540000 0.000000 325.205000 0.630000 ;
      RECT 321.455000 0.000000 323.120000 0.630000 ;
      RECT 319.370000 0.000000 321.035000 0.630000 ;
      RECT 317.280000 0.000000 318.950000 0.630000 ;
      RECT 315.195000 0.000000 316.860000 0.630000 ;
      RECT 313.110000 0.000000 314.775000 0.630000 ;
      RECT 311.025000 0.000000 312.690000 0.630000 ;
      RECT 308.940000 0.000000 310.605000 0.630000 ;
      RECT 306.850000 0.000000 308.520000 0.630000 ;
      RECT 304.765000 0.000000 306.430000 0.630000 ;
      RECT 302.680000 0.000000 304.345000 0.630000 ;
      RECT 300.595000 0.000000 302.260000 0.630000 ;
      RECT 298.510000 0.000000 300.175000 0.630000 ;
      RECT 296.420000 0.000000 298.090000 0.630000 ;
      RECT 294.335000 0.000000 296.000000 0.630000 ;
      RECT 292.250000 0.000000 293.915000 0.630000 ;
      RECT 290.165000 0.000000 291.830000 0.630000 ;
      RECT 288.080000 0.000000 289.745000 0.630000 ;
      RECT 285.990000 0.000000 287.660000 0.630000 ;
      RECT 283.905000 0.000000 285.570000 0.630000 ;
      RECT 281.820000 0.000000 283.485000 0.630000 ;
      RECT 279.735000 0.000000 281.400000 0.630000 ;
      RECT 277.650000 0.000000 279.315000 0.630000 ;
      RECT 275.560000 0.000000 277.230000 0.630000 ;
      RECT 273.475000 0.000000 275.140000 0.630000 ;
      RECT 271.390000 0.000000 273.055000 0.630000 ;
      RECT 269.305000 0.000000 270.970000 0.630000 ;
      RECT 267.220000 0.000000 268.885000 0.630000 ;
      RECT 265.130000 0.000000 266.800000 0.630000 ;
      RECT 263.045000 0.000000 264.710000 0.630000 ;
      RECT 260.960000 0.000000 262.625000 0.630000 ;
      RECT 258.875000 0.000000 260.540000 0.630000 ;
      RECT 256.790000 0.000000 258.455000 0.630000 ;
      RECT 254.700000 0.000000 256.370000 0.630000 ;
      RECT 252.615000 0.000000 254.280000 0.630000 ;
      RECT 250.530000 0.000000 252.195000 0.630000 ;
      RECT 248.445000 0.000000 250.110000 0.630000 ;
      RECT 246.360000 0.000000 248.025000 0.630000 ;
      RECT 244.270000 0.000000 245.940000 0.630000 ;
      RECT 242.185000 0.000000 243.850000 0.630000 ;
      RECT 240.100000 0.000000 241.765000 0.630000 ;
      RECT 238.015000 0.000000 239.680000 0.630000 ;
      RECT 235.930000 0.000000 237.595000 0.630000 ;
      RECT 233.840000 0.000000 235.510000 0.630000 ;
      RECT 231.755000 0.000000 233.420000 0.630000 ;
      RECT 229.670000 0.000000 231.335000 0.630000 ;
      RECT 227.585000 0.000000 229.250000 0.630000 ;
      RECT 225.500000 0.000000 227.165000 0.630000 ;
      RECT 223.410000 0.000000 225.080000 0.630000 ;
      RECT 221.325000 0.000000 222.990000 0.630000 ;
      RECT 219.240000 0.000000 220.905000 0.630000 ;
      RECT 217.155000 0.000000 218.820000 0.630000 ;
      RECT 215.070000 0.000000 216.735000 0.630000 ;
      RECT 212.980000 0.000000 214.650000 0.630000 ;
      RECT 210.895000 0.000000 212.560000 0.630000 ;
      RECT 208.810000 0.000000 210.475000 0.630000 ;
      RECT 206.725000 0.000000 208.390000 0.630000 ;
      RECT 204.640000 0.000000 206.305000 0.630000 ;
      RECT 202.550000 0.000000 204.220000 0.630000 ;
      RECT 200.465000 0.000000 202.130000 0.630000 ;
      RECT 198.380000 0.000000 200.045000 0.630000 ;
      RECT 196.295000 0.000000 197.960000 0.630000 ;
      RECT 194.210000 0.000000 195.875000 0.630000 ;
      RECT 192.120000 0.000000 193.790000 0.630000 ;
      RECT 190.035000 0.000000 191.700000 0.630000 ;
      RECT 187.950000 0.000000 189.615000 0.630000 ;
      RECT 185.865000 0.000000 187.530000 0.630000 ;
      RECT 183.780000 0.000000 185.445000 0.630000 ;
      RECT 181.690000 0.000000 183.360000 0.630000 ;
      RECT 179.605000 0.000000 181.270000 0.630000 ;
      RECT 177.520000 0.000000 179.185000 0.630000 ;
      RECT 175.435000 0.000000 177.100000 0.630000 ;
      RECT 173.350000 0.000000 175.015000 0.630000 ;
      RECT 171.260000 0.000000 172.930000 0.630000 ;
      RECT 169.175000 0.000000 170.840000 0.630000 ;
      RECT 167.090000 0.000000 168.755000 0.630000 ;
      RECT 165.005000 0.000000 166.670000 0.630000 ;
      RECT 162.920000 0.000000 164.585000 0.630000 ;
      RECT 160.830000 0.000000 162.500000 0.630000 ;
      RECT 158.745000 0.000000 160.410000 0.630000 ;
      RECT 156.660000 0.000000 158.325000 0.630000 ;
      RECT 154.575000 0.000000 156.240000 0.630000 ;
      RECT 152.490000 0.000000 154.155000 0.630000 ;
      RECT 150.400000 0.000000 152.070000 0.630000 ;
      RECT 148.315000 0.000000 149.980000 0.630000 ;
      RECT 146.230000 0.000000 147.895000 0.630000 ;
      RECT 144.145000 0.000000 145.810000 0.630000 ;
      RECT 142.060000 0.000000 143.725000 0.630000 ;
      RECT 139.970000 0.000000 141.640000 0.630000 ;
      RECT 137.885000 0.000000 139.550000 0.630000 ;
      RECT 135.800000 0.000000 137.465000 0.630000 ;
      RECT 133.715000 0.000000 135.380000 0.630000 ;
      RECT 131.630000 0.000000 133.295000 0.630000 ;
      RECT 129.540000 0.000000 131.210000 0.630000 ;
      RECT 127.455000 0.000000 129.120000 0.630000 ;
      RECT 125.370000 0.000000 127.035000 0.630000 ;
      RECT 123.285000 0.000000 124.950000 0.630000 ;
      RECT 121.200000 0.000000 122.865000 0.630000 ;
      RECT 119.110000 0.000000 120.780000 0.630000 ;
      RECT 117.025000 0.000000 118.690000 0.630000 ;
      RECT 114.940000 0.000000 116.605000 0.630000 ;
      RECT 112.855000 0.000000 114.520000 0.630000 ;
      RECT 110.770000 0.000000 112.435000 0.630000 ;
      RECT 108.680000 0.000000 110.350000 0.630000 ;
      RECT 106.595000 0.000000 108.260000 0.630000 ;
      RECT 104.510000 0.000000 106.175000 0.630000 ;
      RECT 102.425000 0.000000 104.090000 0.630000 ;
      RECT 100.340000 0.000000 102.005000 0.630000 ;
      RECT 98.250000 0.000000 99.920000 0.630000 ;
      RECT 96.165000 0.000000 97.830000 0.630000 ;
      RECT 94.080000 0.000000 95.745000 0.630000 ;
      RECT 91.995000 0.000000 93.660000 0.630000 ;
      RECT 89.910000 0.000000 91.575000 0.630000 ;
      RECT 87.820000 0.000000 89.490000 0.630000 ;
      RECT 85.735000 0.000000 87.400000 0.630000 ;
      RECT 83.650000 0.000000 85.315000 0.630000 ;
      RECT 81.565000 0.000000 83.230000 0.630000 ;
      RECT 79.480000 0.000000 81.145000 0.630000 ;
      RECT 77.390000 0.000000 79.060000 0.630000 ;
      RECT 75.305000 0.000000 76.970000 0.630000 ;
      RECT 73.220000 0.000000 74.885000 0.630000 ;
      RECT 71.135000 0.000000 72.800000 0.630000 ;
      RECT 69.050000 0.000000 70.715000 0.630000 ;
      RECT 66.960000 0.000000 68.630000 0.630000 ;
      RECT 64.875000 0.000000 66.540000 0.630000 ;
      RECT 62.790000 0.000000 64.455000 0.630000 ;
      RECT 60.705000 0.000000 62.370000 0.630000 ;
      RECT 58.620000 0.000000 60.285000 0.630000 ;
      RECT 56.530000 0.000000 58.200000 0.630000 ;
      RECT 54.445000 0.000000 56.110000 0.630000 ;
      RECT 52.360000 0.000000 54.025000 0.630000 ;
      RECT 50.275000 0.000000 51.940000 0.630000 ;
      RECT 48.190000 0.000000 49.855000 0.630000 ;
      RECT 46.100000 0.000000 47.770000 0.630000 ;
      RECT 44.015000 0.000000 45.680000 0.630000 ;
      RECT 41.930000 0.000000 43.595000 0.630000 ;
      RECT 39.845000 0.000000 41.510000 0.630000 ;
      RECT 37.760000 0.000000 39.425000 0.630000 ;
      RECT 35.670000 0.000000 37.340000 0.630000 ;
      RECT 33.585000 0.000000 35.250000 0.630000 ;
      RECT 31.500000 0.000000 33.165000 0.630000 ;
      RECT 29.415000 0.000000 31.080000 0.630000 ;
      RECT 27.330000 0.000000 28.995000 0.630000 ;
      RECT 25.240000 0.000000 26.910000 0.630000 ;
      RECT 23.155000 0.000000 24.820000 0.630000 ;
      RECT 21.070000 0.000000 22.735000 0.630000 ;
      RECT 18.985000 0.000000 20.650000 0.630000 ;
      RECT 16.900000 0.000000 18.565000 0.630000 ;
      RECT 14.810000 0.000000 16.480000 0.630000 ;
      RECT 12.725000 0.000000 14.390000 0.630000 ;
      RECT 10.640000 0.000000 12.305000 0.630000 ;
      RECT 8.555000 0.000000 10.220000 0.630000 ;
      RECT 6.470000 0.000000 8.135000 0.630000 ;
      RECT 4.380000 0.000000 6.050000 0.630000 ;
      RECT 2.295000 0.000000 3.960000 0.630000 ;
      RECT 0.000000 0.000000 1.875000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 1015.150000 1020.280000 1019.660000 ;
      RECT 1.100000 1014.540000 1020.280000 1015.150000 ;
      RECT 1.100000 1014.250000 1019.180000 1014.540000 ;
      RECT 0.000000 1013.640000 1019.180000 1014.250000 ;
      RECT 0.000000 996.930000 1020.280000 1013.640000 ;
      RECT 0.000000 996.030000 1019.180000 996.930000 ;
      RECT 0.000000 995.210000 1020.280000 996.030000 ;
      RECT 1.100000 994.310000 1020.280000 995.210000 ;
      RECT 0.000000 973.760000 1020.280000 994.310000 ;
      RECT 0.000000 972.860000 1019.180000 973.760000 ;
      RECT 0.000000 970.340000 1020.280000 972.860000 ;
      RECT 1.100000 969.440000 1020.280000 970.340000 ;
      RECT 0.000000 950.585000 1020.280000 969.440000 ;
      RECT 0.000000 949.685000 1019.180000 950.585000 ;
      RECT 0.000000 945.470000 1020.280000 949.685000 ;
      RECT 1.100000 944.570000 1020.280000 945.470000 ;
      RECT 0.000000 927.410000 1020.280000 944.570000 ;
      RECT 0.000000 926.510000 1019.180000 927.410000 ;
      RECT 0.000000 920.605000 1020.280000 926.510000 ;
      RECT 1.100000 919.705000 1020.280000 920.605000 ;
      RECT 0.000000 904.235000 1020.280000 919.705000 ;
      RECT 0.000000 903.335000 1019.180000 904.235000 ;
      RECT 0.000000 895.735000 1020.280000 903.335000 ;
      RECT 1.100000 894.835000 1020.280000 895.735000 ;
      RECT 0.000000 881.060000 1020.280000 894.835000 ;
      RECT 0.000000 880.160000 1019.180000 881.060000 ;
      RECT 0.000000 870.865000 1020.280000 880.160000 ;
      RECT 1.100000 869.965000 1020.280000 870.865000 ;
      RECT 0.000000 857.890000 1020.280000 869.965000 ;
      RECT 0.000000 856.990000 1019.180000 857.890000 ;
      RECT 0.000000 845.995000 1020.280000 856.990000 ;
      RECT 1.100000 845.095000 1020.280000 845.995000 ;
      RECT 0.000000 834.715000 1020.280000 845.095000 ;
      RECT 0.000000 833.815000 1019.180000 834.715000 ;
      RECT 0.000000 821.125000 1020.280000 833.815000 ;
      RECT 1.100000 820.225000 1020.280000 821.125000 ;
      RECT 0.000000 811.540000 1020.280000 820.225000 ;
      RECT 0.000000 810.640000 1019.180000 811.540000 ;
      RECT 0.000000 796.260000 1020.280000 810.640000 ;
      RECT 1.100000 795.360000 1020.280000 796.260000 ;
      RECT 0.000000 788.365000 1020.280000 795.360000 ;
      RECT 0.000000 787.465000 1019.180000 788.365000 ;
      RECT 0.000000 771.390000 1020.280000 787.465000 ;
      RECT 1.100000 770.490000 1020.280000 771.390000 ;
      RECT 0.000000 765.190000 1020.280000 770.490000 ;
      RECT 0.000000 764.290000 1019.180000 765.190000 ;
      RECT 0.000000 746.520000 1020.280000 764.290000 ;
      RECT 1.100000 745.620000 1020.280000 746.520000 ;
      RECT 0.000000 742.020000 1020.280000 745.620000 ;
      RECT 0.000000 741.120000 1019.180000 742.020000 ;
      RECT 0.000000 721.650000 1020.280000 741.120000 ;
      RECT 1.100000 720.750000 1020.280000 721.650000 ;
      RECT 0.000000 718.845000 1020.280000 720.750000 ;
      RECT 0.000000 717.945000 1019.180000 718.845000 ;
      RECT 0.000000 696.780000 1020.280000 717.945000 ;
      RECT 1.100000 695.880000 1020.280000 696.780000 ;
      RECT 0.000000 695.670000 1020.280000 695.880000 ;
      RECT 0.000000 694.770000 1019.180000 695.670000 ;
      RECT 0.000000 672.495000 1020.280000 694.770000 ;
      RECT 0.000000 671.915000 1019.180000 672.495000 ;
      RECT 1.100000 671.595000 1019.180000 671.915000 ;
      RECT 1.100000 671.015000 1020.280000 671.595000 ;
      RECT 0.000000 649.320000 1020.280000 671.015000 ;
      RECT 0.000000 648.420000 1019.180000 649.320000 ;
      RECT 0.000000 647.045000 1020.280000 648.420000 ;
      RECT 1.100000 646.145000 1020.280000 647.045000 ;
      RECT 0.000000 626.150000 1020.280000 646.145000 ;
      RECT 0.000000 625.250000 1019.180000 626.150000 ;
      RECT 0.000000 622.175000 1020.280000 625.250000 ;
      RECT 1.100000 621.275000 1020.280000 622.175000 ;
      RECT 0.000000 602.975000 1020.280000 621.275000 ;
      RECT 0.000000 602.075000 1019.180000 602.975000 ;
      RECT 0.000000 597.305000 1020.280000 602.075000 ;
      RECT 1.100000 596.405000 1020.280000 597.305000 ;
      RECT 0.000000 579.800000 1020.280000 596.405000 ;
      RECT 0.000000 578.900000 1019.180000 579.800000 ;
      RECT 0.000000 572.435000 1020.280000 578.900000 ;
      RECT 1.100000 571.535000 1020.280000 572.435000 ;
      RECT 0.000000 556.625000 1020.280000 571.535000 ;
      RECT 0.000000 555.725000 1019.180000 556.625000 ;
      RECT 0.000000 547.570000 1020.280000 555.725000 ;
      RECT 1.100000 546.670000 1020.280000 547.570000 ;
      RECT 0.000000 533.450000 1020.280000 546.670000 ;
      RECT 0.000000 532.550000 1019.180000 533.450000 ;
      RECT 0.000000 522.700000 1020.280000 532.550000 ;
      RECT 1.100000 521.800000 1020.280000 522.700000 ;
      RECT 0.000000 510.280000 1020.280000 521.800000 ;
      RECT 0.000000 509.380000 1019.180000 510.280000 ;
      RECT 0.000000 497.830000 1020.280000 509.380000 ;
      RECT 1.100000 496.930000 1020.280000 497.830000 ;
      RECT 0.000000 487.105000 1020.280000 496.930000 ;
      RECT 0.000000 486.205000 1019.180000 487.105000 ;
      RECT 0.000000 472.960000 1020.280000 486.205000 ;
      RECT 1.100000 472.060000 1020.280000 472.960000 ;
      RECT 0.000000 463.930000 1020.280000 472.060000 ;
      RECT 0.000000 463.030000 1019.180000 463.930000 ;
      RECT 0.000000 448.090000 1020.280000 463.030000 ;
      RECT 1.100000 447.190000 1020.280000 448.090000 ;
      RECT 0.000000 440.755000 1020.280000 447.190000 ;
      RECT 0.000000 439.855000 1019.180000 440.755000 ;
      RECT 0.000000 423.225000 1020.280000 439.855000 ;
      RECT 1.100000 422.325000 1020.280000 423.225000 ;
      RECT 0.000000 417.580000 1020.280000 422.325000 ;
      RECT 0.000000 416.680000 1019.180000 417.580000 ;
      RECT 0.000000 398.355000 1020.280000 416.680000 ;
      RECT 1.100000 397.455000 1020.280000 398.355000 ;
      RECT 0.000000 394.410000 1020.280000 397.455000 ;
      RECT 0.000000 393.510000 1019.180000 394.410000 ;
      RECT 0.000000 373.485000 1020.280000 393.510000 ;
      RECT 1.100000 372.585000 1020.280000 373.485000 ;
      RECT 0.000000 371.235000 1020.280000 372.585000 ;
      RECT 0.000000 370.335000 1019.180000 371.235000 ;
      RECT 0.000000 348.615000 1020.280000 370.335000 ;
      RECT 1.100000 348.060000 1020.280000 348.615000 ;
      RECT 1.100000 347.715000 1019.180000 348.060000 ;
      RECT 0.000000 347.160000 1019.180000 347.715000 ;
      RECT 0.000000 324.885000 1020.280000 347.160000 ;
      RECT 0.000000 323.985000 1019.180000 324.885000 ;
      RECT 0.000000 323.745000 1020.280000 323.985000 ;
      RECT 1.100000 322.845000 1020.280000 323.745000 ;
      RECT 0.000000 301.710000 1020.280000 322.845000 ;
      RECT 0.000000 300.810000 1019.180000 301.710000 ;
      RECT 0.000000 298.880000 1020.280000 300.810000 ;
      RECT 1.100000 297.980000 1020.280000 298.880000 ;
      RECT 0.000000 278.540000 1020.280000 297.980000 ;
      RECT 0.000000 277.640000 1019.180000 278.540000 ;
      RECT 0.000000 274.010000 1020.280000 277.640000 ;
      RECT 1.100000 273.110000 1020.280000 274.010000 ;
      RECT 0.000000 255.365000 1020.280000 273.110000 ;
      RECT 0.000000 254.465000 1019.180000 255.365000 ;
      RECT 0.000000 249.140000 1020.280000 254.465000 ;
      RECT 1.100000 248.240000 1020.280000 249.140000 ;
      RECT 0.000000 232.190000 1020.280000 248.240000 ;
      RECT 0.000000 231.290000 1019.180000 232.190000 ;
      RECT 0.000000 224.270000 1020.280000 231.290000 ;
      RECT 1.100000 223.370000 1020.280000 224.270000 ;
      RECT 0.000000 209.015000 1020.280000 223.370000 ;
      RECT 0.000000 208.115000 1019.180000 209.015000 ;
      RECT 0.000000 199.400000 1020.280000 208.115000 ;
      RECT 1.100000 198.500000 1020.280000 199.400000 ;
      RECT 0.000000 185.840000 1020.280000 198.500000 ;
      RECT 0.000000 184.940000 1019.180000 185.840000 ;
      RECT 0.000000 174.535000 1020.280000 184.940000 ;
      RECT 1.100000 173.635000 1020.280000 174.535000 ;
      RECT 0.000000 162.670000 1020.280000 173.635000 ;
      RECT 0.000000 161.770000 1019.180000 162.670000 ;
      RECT 0.000000 149.665000 1020.280000 161.770000 ;
      RECT 1.100000 148.765000 1020.280000 149.665000 ;
      RECT 0.000000 139.495000 1020.280000 148.765000 ;
      RECT 0.000000 138.595000 1019.180000 139.495000 ;
      RECT 0.000000 124.795000 1020.280000 138.595000 ;
      RECT 1.100000 123.895000 1020.280000 124.795000 ;
      RECT 0.000000 116.320000 1020.280000 123.895000 ;
      RECT 0.000000 115.420000 1019.180000 116.320000 ;
      RECT 0.000000 99.925000 1020.280000 115.420000 ;
      RECT 1.100000 99.025000 1020.280000 99.925000 ;
      RECT 0.000000 93.145000 1020.280000 99.025000 ;
      RECT 0.000000 92.245000 1019.180000 93.145000 ;
      RECT 0.000000 75.055000 1020.280000 92.245000 ;
      RECT 1.100000 74.155000 1020.280000 75.055000 ;
      RECT 0.000000 69.970000 1020.280000 74.155000 ;
      RECT 0.000000 69.070000 1019.180000 69.970000 ;
      RECT 0.000000 50.190000 1020.280000 69.070000 ;
      RECT 1.100000 49.290000 1020.280000 50.190000 ;
      RECT 0.000000 46.800000 1020.280000 49.290000 ;
      RECT 0.000000 45.900000 1019.180000 46.800000 ;
      RECT 0.000000 25.320000 1020.280000 45.900000 ;
      RECT 1.100000 24.420000 1020.280000 25.320000 ;
      RECT 0.000000 23.625000 1020.280000 24.420000 ;
      RECT 0.000000 22.725000 1019.180000 23.625000 ;
      RECT 0.000000 20.850000 1020.280000 22.725000 ;
      RECT 1.100000 19.950000 1020.280000 20.850000 ;
      RECT 0.000000 10.480000 1020.280000 19.950000 ;
      RECT 1.100000 9.580000 1020.280000 10.480000 ;
      RECT 0.000000 4.990000 1020.280000 9.580000 ;
      RECT 0.000000 4.090000 1019.180000 4.990000 ;
      RECT 0.000000 1.330000 1020.280000 4.090000 ;
      RECT 1.100000 1.100000 1020.280000 1.330000 ;
      RECT 1.100000 0.430000 4.380000 1.100000 ;
      RECT 5.280000 0.000000 1020.280000 1.100000 ;
      RECT 0.000000 0.000000 4.380000 0.430000 ;
    LAYER met4 ;
      RECT 0.000000 1017.180000 1020.280000 1019.660000 ;
      RECT 4.360000 1013.180000 1015.920000 1017.180000 ;
      RECT 1014.520000 5.630000 1015.920000 1013.180000 ;
      RECT 8.360000 5.630000 1011.920000 1013.180000 ;
      RECT 4.360000 5.630000 5.760000 1013.180000 ;
      RECT 1018.520000 1.630000 1020.280000 1017.180000 ;
      RECT 4.360000 1.630000 1015.920000 5.630000 ;
      RECT 0.000000 1.630000 1.760000 1017.180000 ;
      RECT 0.000000 0.000000 1020.280000 1.630000 ;
  END
END user_proj_example

END LIBRARY
